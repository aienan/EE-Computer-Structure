`timescale 1ns/1ns

module tb_SimpleMIPS;
    reg clk, rstn, im_write;
    reg [31:0] im_addr;
    reg [31:0] im_wdata;
        
    SimpleMIPS a_0(.clk(clk), .rstn(rstn), .im_write(im_write), .im_addr(im_addr), .im_wdata(im_wdata));
    
    initial begin
       clk <= 1;
	    forever #5 clk <= ~clk;
    end
    
    initial begin
       im_write <= 1;
       rstn <= 1;
              
       #20
       im_addr <= 1;
       im_wdata <= 32'b 000100_00000_00001_0000_0000_1011_0010;      // addi $s1, $s0, 178
       #20
       im_addr <= 2;
       im_wdata <= 32'b 000100_00000_00010_0000_0000_0000_1100;      // addi $s2, $s0, 12
       #20
       im_addr <= 3;
       im_wdata <= 32'b 000011_00001_00010_0001_1000_0000_0000;      // add $s3, $s1, $s2
       #20
       im_addr <= 4;
       im_wdata <= 32'b 000101_00001_00010_0010_0000_0000_0000;      // sub $s4, $s1, $s2
       #20
       im_addr <= 5;
       im_wdata <= 32'b 000100_00001_00101_0000_0000_0000_0000;      // addi $s5, $s1, 0
       #20
       im_addr <= 6;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 7;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 8;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 9;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 10;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 11;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 12;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 13;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 14;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 15;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 16;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 17;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 18;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 19;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 20;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 21;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 22;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 23;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 24;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 25;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 26;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 27;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 28;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 29;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 30;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 31;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 32;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 33;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 34;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 35;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 36;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
       #20
       im_addr <= 37;
       im_wdata <= 32'b 000110_00101_00010_0010_1000_0000_0000;      // div $s5, $s5, $s2
              
        
       #20
       im_write <= 0;
       
       #20
       rstn <= 0;
        
        
        
        
    end
    
endmodule